    <svg
              aria-hidden="true"
              focusable="false"
              data-prefix="far"
              data-icon="arrow-turn-up"
              class="svg-inline--fa fa-arrow-turn-up fa-flip-horizontal"
              role="img"
              xmlns="http://www.w3.org/2000/svg"
              viewBox="0 0 384 512"
            >
              <path
                fill="currentColor"
                d="M24 464c-13.3 0-24 10.7-24 24s10.7 24 24 24l104 0c48.6 0 88-39.4 88-88l0-342.1 87 87c9.4 9.4 24.6 9.4 33.9 0s9.4-24.6 0-33.9L209 7c-9.4-9.4-24.6-9.4-33.9 0L47 135c-9.4 9.4-9.4 24.6 0 33.9s24.6 9.4 33.9 0l87-87L168 424c0 22.1-17.9 40-40 40L24 464z"
              ></path>
            </svg>